`timescale 1ns/1ps

module top (
    input wire clk
    );


    always_ff @(posedge clk) begin
        
    end
endmodule
