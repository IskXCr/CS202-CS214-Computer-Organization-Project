`timescale 1ns/1ps

module beeper(

    );
    
endmodule