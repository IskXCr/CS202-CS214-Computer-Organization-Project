`timescale 1ns/1ps

module cpu_sim();
    
    always begin
        
    end
endmodule