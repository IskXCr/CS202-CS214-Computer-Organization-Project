`timescale 1ns/1ps

module top (
    input  wire clk,
    input  wire rst
    );

    wire cpu_clk;
    
    wire mem_write;
    wire [31:0] instr_addr, instr, mem_addr, write_data;
    reg  [31:0] read_data;
    
//    clk_wiz_0 clk_gen(.clk_in1(clk),
//                      .clk_out1(cpu_clk));
    assign cpu_clk = clk;
                          
    CPU cpu_inst(.clk(cpu_clk),
                 .rst(rst),
                 .instr_addr(instr_addr),
                 .instr(instr),
                 .mem_write(mem_write),
                 .mem_addr(mem_addr),
                 .write_data(write_data),
                 .read_data(read_data));
    
    // set instruction memory
    wire [31:0] true_instr_addr;
    
    assign true_instr_addr = $signed(instr_addr) - $signed(32'h0040_0000);
                 
    instr_mem instr_memory(.clka(cpu_clk),
                           .addra(true_instr_addr[15:2]),
                           .wea(0),
                           .dina(0),
                           .douta(instr));
    
    // set data memory
    wire is_in_data_seg;
    wire [31:0] data_addr;
    wire data_wea;
    wire data_out;
    
    assign is_in_data_seg = (mem_addr >= 32'h7fff000 && mem_addr <= 32'h7fffeffc);
    assign data_addr = is_in_data_seg ? ($signed(mem_addr) - $signed(32'h1001_0000)) : 32'h00000000;
    assign data_wea = is_in_data_seg && mem_write;
    
    data_mem data_memory(.clka(~cpu_clk),
                         .addra(data_addr[15:2]),
                         .dina(write_data),
                         .douta(data_out),
                         .wea(data_wea));
    
    // set stack memory
    wire is_in_stack_seg;
    wire [31:0] stack_addr;
    wire stack_wea;
    wire stack_out;
    
    assign is_in_stack_seg = (mem_addr >= 32'h7fff000 && mem_addr <= 32'h7fffeffc);
    assign stack_addr = is_in_stack_seg  ? (32'h7fffeffc - mem_addr) : 32'h00000000;
    assign stack_wea = is_in_stack_seg  && mem_write;
    
    stack_mem stack_memory(.clka(~cpu_clk),
                           .addra(stack_addr[15:2]),
                           .dina(write_data),
                           .douta(stack_out),
                           .wea(stack_wea));
    
    
    // set the source of read_data
    wire [1:0] data_dst;
    
    assign data_dst = {is_in_data_seg, is_in_stack_seg};
    
    // adjust read port
    always_comb begin
        casez (data_dst)
            2'b10: read_data = data_out;
            2'b01: read_data = stack_out;
            default: read_data = 32'h00000000;
        endcase
    end
    
endmodule
