`timescale 1ns/1ps

module top (
    input  wire cpu_clk,
    input  wire mem_clk
    );


    always_ff @(posedge clk) begin
        
    end
endmodule
