`timescale 1ns / 1ps

module controller (
    input  wire clk,
    input  wire [31:0] inst
    );


    always_ff @(posedge clk) begin
        
    end
endmodule
