`timescale 1ns/1ps

module inst_fetch (
    input wire clk
    );


    always_ff @(posedge clk) begin
        
    end
endmodule
